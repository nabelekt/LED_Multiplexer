** Profile: "SCHEMATIC1-multiplexer_sim"  [ \\aerobus3\Users6$\tnabelek\My Documents\Development Projects\LED Multiplexer\LED Multiplexer-PSpiceFiles\SCHEMATIC1\multiplexer_sim.sim ] 

** Creating circuit file "multiplexer_sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
