** Profile: "SCHEMATIC1-Potentiometer_Sweep"  [ C:\Users\Thomas Nabelek\Desktop\LED_Multiplexer\stage_2\led multiplexer-pspicefiles\schematic1\potentiometer_sweep.sim ] 

** Creating circuit file "Potentiometer_Sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN PARAM OHM 30 200 1 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
