** Profile: "SCHEMATIC1-transistor_r_sweep"  [ \\aerobus3\Users6$\tnabelek\My Documents\Development Projects\LED_Multiplexer\stage_2\LED Multiplexer-PSpiceFiles\SCHEMATIC1\transistor_r_sweep.sim ] 

** Creating circuit file "transistor_r_sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\tnabelek\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN PARAM TRANSISTOR_R 1 50000 20 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
